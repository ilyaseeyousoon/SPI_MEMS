module centroids (input clk_200MHz_i,
					input rdempty,
					input start_treatment,
					input reset,
					input [20:0] window_input,
					input [29:0] numerator,
					output clken,
					output read_fifo,
					output aclr_fifo,
					output [20:0] denominator );
					
					
					
					
endmodule