library verilog;
use verilog.vl_types.all;
entity clk_to_ADC_tb is
end clk_to_ADC_tb;
