library verilog;
use verilog.vl_types.all;
entity top_file_vlg_tst is
end top_file_vlg_tst;
