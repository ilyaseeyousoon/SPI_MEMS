module counter_reset_diods  (input clk_5MHz_i,output [15:0] n );

endmodule