library verilog;
use verilog.vl_types.all;
entity firsttry_tb is
end firsttry_tb;
