// megafunction wizard: %LPM_DIVIDE%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_DIVIDE 

// ============================================================
// File Name: div_first.v
// Megafunction Name(s):
// 			LPM_DIVIDE
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 14.0.0 Build 200 06/17/2014 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, the Altera Quartus II License Agreement,
//the Altera MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Altera and sold by Altera or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.

module div_first (
	clken,
	clock,
	denom,
	numer,
	quotient,
	remain);

	input	  clken;
	input	  clock;
	input	[26:0]  denom;
	input	[39:0]  numer;
	output	[39:0]  quotient;
	output	[26:0]  remain;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE"
// Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "-1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "1"
// Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_HINT STRING "LPM_REMAINDERPOSITIVE=TRUE"
// Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "40"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
// Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "27"
// Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "40"
// Retrieval info: USED_PORT: clken 0 0 0 0 INPUT NODEFVAL "clken"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: denom 0 0 27 0 INPUT NODEFVAL "denom[26..0]"
// Retrieval info: USED_PORT: numer 0 0 40 0 INPUT NODEFVAL "numer[39..0]"
// Retrieval info: USED_PORT: quotient 0 0 40 0 OUTPUT NODEFVAL "quotient[39..0]"
// Retrieval info: USED_PORT: remain 0 0 27 0 OUTPUT NODEFVAL "remain[26..0]"
// Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @denom 0 0 27 0 denom 0 0 27 0
// Retrieval info: CONNECT: @numer 0 0 40 0 numer 0 0 40 0
// Retrieval info: CONNECT: quotient 0 0 40 0 @quotient 0 0 40 0
// Retrieval info: CONNECT: remain 0 0 27 0 @remain 0 0 27 0
// Retrieval info: GEN_FILE: TYPE_NORMAL div_first.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_first.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_first.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_first.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_first_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_first_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
