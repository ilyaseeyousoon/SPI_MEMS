module concatenation   (			
										input clk_200MHz_i,
										input wful,
										input remp,
										input [39:0] quot,
										input [7:0] rem,
										output  rdreq,
										output centroid_out );
										


										
assign rdreq=0;										
endmodule