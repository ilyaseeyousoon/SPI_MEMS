module filtered_adc_data_to_fifo  (input clk_5MHz_i,output [15:0] n );

endmodule