module wait_signals_AD_sp_and_AD_trig  (input clk_5MHz_i,output [15:0] n );

endmodule